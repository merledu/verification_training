class porsche extends car;
  function new(string c="BLACK");
    $display("In Porsche");
  endfunction  
endclass
Porsche p_h=new();