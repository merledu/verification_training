interface intf();

logic [2:0] opA_i;
logic [2:0] opB_i;
modport intf_tb(output opA_i,opB_i);  

endinterface
