class cat extends animal;
  function new();
    weight = 5;
    color = "grey";
  endfunction
endclass