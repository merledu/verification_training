class Vector #(parameter SIZE = 32);
  bit [SIZE-1:0] data;
endclass