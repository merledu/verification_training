package pkg;
  typedef class car;
  typedef class porsche;
  
  `include "car.svh"
  `include "porsche.svh"
endpackage