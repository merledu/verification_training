package pkg;
  // Classes are defined to be used in the virtual interface
  typedef class Driver;
  `include "driver.svh"
endpackage