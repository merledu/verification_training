package pkg;
  typedef class transaction;
  typedef class BadTr;

  `include "transaction.svh"
  `include "BadTr.svh"
endpackage