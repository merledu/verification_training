class animal;
  int weight;
  protected string color;
  local int age;
endclass