class car;
  string color;
  function new(string c="BLACK");
    color = c;
    $display("In Car");
  endfunction
endclass            