module test();
  
  typedef class Animal;
  typedef class Mouth;
  
  Animal a_h;

  class Animal;
    Mouth a_h;

  endclass
endmodule