package pkg;
  typedef class Animal;
  typedef class Cat;
  `include "Animal_class.svh"
  `include "Cat_class.svh"
endpackage