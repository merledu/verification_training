package pkg;
  typedef class animal;
  typedef class cat;

  `include "animal.svh"
  `include "cat.svh"
endpackage