package pkg;
  // Classes are defined to be used
  typedef class Driver;
  `include "driver.svh"
endpackage