/////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:        MICRO-ELECTRONICS RESEARCH LABORATORY                                               //
//                                                                                                     //
// Engineers:      Wishah Naseer - Verification	Engineer                                               //
//                                                                                                     //
// Additional contributions by:                                                                        //
//                                                                                                     //
// Create Date:    20-MARCH-2022                                                                       //
// Design Name:    SV OOP Practice                                                                     //
// Module Name:    Example 06.sv                                                                       //
// Project Name:   SV OOP Training                                                                     //
// Language:       SystemVerilog - UVM                                                                 //
//                                                                                                     //
// Description:                                                                                        //
//     - This code helps to understand how multiple handles can point to a single object.  ....	       //
//                                                                                                     //
//                                                                                                     //
// Revision Date:                                                                                      //
//                                                                                                     //
/////////////////////////////////////////////////////////////////////////////////////////////////////////

module top();  
	class Animal;  //class declaration
    //property 
    int age;
    string name;

    //constructor method
    function new(string name, int age); //configurable constructor with same local variables as property
      this.age = age;
      this.name = name;
    endfunction

    //another method
    function void print();
    $display("Animal : '%s' age = a0d", name, age);
    endfunction
    
  endclass : Animal

//multiple handles can point to same object

Animal a1_h;
Animal a2_h;

initial begin
  a1_h = new(.name("Puppy"), .age(5));
  a2_h = a1_h;
end
endmodule
