class usb_monitor;
  
endclass