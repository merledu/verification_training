package pkg;
  typedef class Transaction;
  typedef class BadTr;
  `include "Transaction.svh"
  `include "BadTr.svh"
endpackage