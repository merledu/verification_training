module usb_pkg;

typedef class usb_driver;
typedef class usb_monitor;


`include "usb_driver.svh"
`include "usb_monitor.svh"

endmodule