package pkg;
  typedef class Transaction;
  typedef class BadTr;
  typedef class Generator;
  typedef class BaseTest;
  typedef class BadTest;
  
  
  `include "Transaction.svh"
  `include "BadTr.svh"
  `include "Generator.svh"
  `include "BaseTest.svh"
  `include "BadTest.svh"
endpackage