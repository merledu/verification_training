class usb_driver;
  
endclass