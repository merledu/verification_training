class BaseTest;
  Generator gen_h;

  function new();
    gen_h = new();
  endfunction

  task run();
    gen_h.run();
  endtask

endclass
