module test();
  import usb_pkg::;
  
  usb_driver drv;
  usb_monitor mon;
  
endmodule